netcdf C:/Ethan/code/threddsDev/cdm/src/test/data/dmsp/F14200307192230.n.OIS {
 dimensions:
   numScans = 691;
   numSamplesPerScan = 1465;
 variables:
   int year(numScans=691);
     :long_name = "year at time of scan";
     :units = "year";
   int dayOfYear(numScans=691);
     :long_name = "day of year at time of scan";
     :units = "day of year";
   double secondsOfDay(numScans=691);
     :long_name = "seconds of day at time of scan";
     :units = "seconds of day";
   float time(numScans=691);
     :long_name = "time of scan";
     :units = "seconds since 2003-07-19T22:30:31.371GMT";
     :calculatedVariable = "Using the satellite epoch for each scan.";
     :_CoordinateAxisType = "Time";
   float satEphemLatitude(numScans=691);
     :long_name = "geodetic latitude of the satellite for this scan";
     :units = "degrees_north";
   float satEphemLongitude(numScans=691);
     :long_name = "longitude of the satellite for this scan";
     :units = "degrees_east";
   float satEphemAltitude(numScans=691);
     :long_name = "altitude of the satellite for this scan";
     :units = "kilometers";
   float satEphemHeading(numScans=691);
     :long_name = "heading of the satellite (degrees west of north) for this scan";
     :units = "degrees";
   float scannerOffset(numScans=691);
     :long_name = "scanner offset";
     :units = "radians";
   byte scanDirection(numScans=691);
     :long_name = "scan direction";
     :units = "";
   float solarElevation(numScans=691);
     :long_name = "solar elevation";
     :units = "degrees";
   float solarAzimuth(numScans=691);
     :long_name = "solar azimuth";
     :units = "degrees";
   float lunarElevation(numScans=691);
     :long_name = "lunar elevation";
     :units = "degrees";
   float lunarAzimuth(numScans=691);
     :long_name = "lunar azimuth";
     :units = "degrees";
   float lunarPhase(numScans=691);
     :long_name = "lunar phase";
     :units = "degrees";
   float gainCode(numScans=691);
     :long_name = "gain code";
     :units = "decibels";
   byte gainMode(numScans=691);
     :long_name = "gain mode (0=linear, 1=logrithmic)";
     :units = "";
   byte gainSubMode(numScans=691);
     :long_name = "gain sub-mode";
     :units = "";
   byte hotTCalSegmentID(numScans=691);
     :long_name = "Hot T cal seg ID (0 = right, 1 = left)";
     :units = "";
   byte coldTCalSegmentID(numScans=691);
     :long_name = "Cold T cal seg ID (0 = right, 1 = left)";
     :units = "";
   byte hotTCal(numScans=691);
     :long_name = "Hot T calibration";
     :units = "";
   byte coldTCal(numScans=691);
     :long_name = "Cold T calibration";
     :units = "";
   byte pmtCal(numScans=691);
     :long_name = "Photomultiplier tube calibration";
     :units = "";
   float tChannelGain(numScans=691);
     :long_name = "T channel gain";
     :units = "decibels";
   int visibleScanQualityFlag(numScans=691);
     :long_name = "quality flag for the visible scan";
     :units = "";
   int thermalScanQualityFlag(numScans=691);
     :long_name = "quality flag for the thermal scan";
     :units = "";
   float latitude(numScans=691, numSamplesPerScan=1465);
     :long_name = "latitude of pixel";
     :units = "degrees_north";
     :calculatedVariable = "Using the geometry of the satellite scans and an ellipsoidal earth (a=6378.14km and e=0.0818191830).";
     :_CoordinateAxisType = "Lat";
   float longitude(numScans=691, numSamplesPerScan=1465);
     :long_name = "longitude of pixel";
     :units = "degrees_east";
     :calculatedVariable = "Using the geometry of the satellite scans and an ellipsoidal earth (a=6378.14km and e=0.0818191830).";
     :_CoordinateAxisType = "Lon";
   byte visibleImagery(numScans=691, numSamplesPerScan=1465);
     :long_name = "visible imagery  (6-bit per pixel)";
     :units = "";
     :_CoordinateAxes = "latitude longitude";
     :_unsigned = "true";
     :description = "Visible pixels are relative values ranging from 0 to 63 rather than absolute values in Watts per m^2. Instrumental gain levels are adjusted to maintain constant cloud reference values under varying conditions of solar and lunar illumination. Telescope pixel values are replaced by Photo Multiplier Tube (PMT) values at night. -- From http://dmsp.ngdc.noaa.gov/html/sensors/doc_ols.html";
   byte infraredImagery(numScans=691, numSamplesPerScan=1465);
     :long_name = "infrared imagery (8-bit per pixel)";
     :units = "kelvin";
     :_CoordinateAxes = "latitude longitude";
     :_unsigned = "false";
     :scale_factor = 0.47058824f; // float
     :add_offset = 190.0f; // float
     :description = "Infrared pixel values correspond to a temperature range of 190 to 310 Kelvins in 256 equally spaced steps. Onboard calibration is performed during each scan. -- From http://dmsp.ngdc.noaa.gov/html/sensors/doc_ols.html";

 :fileId = "/dmsp/moby-1-3/subscriptions/IBAMA/1353226646955.tmp";
 :datasetId = "DMSP F14 OLS LS & TS";
 :suborbitHistory = "F14200307192230.OIS (1,691)";
 :processingSystem = "v2.1b";
 :processingDate = "2003-07-19T19:33:23.000GMT";
 :spacecraftId = "F14";
 :noradId = "24753";
 :startDate = "2003-07-19T22:30:31.371GMT";
 :endDate = "2003-07-19T22:35:21.836GMT";
 :startDateLocal = "start date local";
 :startTimeLocal = "start time local";
 :startLatitude = 0.0; // double
 :startLongitude = 320.54; // double
 :endLatitude = 16.99; // double
 :endLongitude = 316.69; // double
 :startSubsolarCoords = "20.87 202.37";
 :endSubsolarCoords = "20.87 201.16";
 :startLunarCoords = "UNKNOWN";
 :endLunarCoords = "UNKNOWN";
 :ascendingNode = 320.55; // double
 :nodeHeading = 8.64; // double
 :nominalResolution = "2.7 km";
 :bandsPerScanline = 2; // int
 :bytesPerSample = 1; // int
 :byteOffsetBand1 = 96; // int
 :byteOffsetBand2 = 1568; // int
 :band1 = "OLS Visible .4-1.1um";
 :band2 = "OLS Thermal 10.5-12.6um";
 :bandOrganization = "band interleaved by line";
 :thermalOffset = "190.00 K";
 :thermalScale = "0.47";
 :percentDaylight = 0.0; // double
 :percentFullMoon = 57.8; // double
 :percentTerminatorEvident = 0.0; // double
 :qcFlags = "0=not QC'ed  1=artificial  2=bad vis";
 :title = "NGDC archived DMSP F14 OLS LS & TS data with start time 2003-07-19T22:30:31.371GMT";
 :Convention = "_Coordinates";
 :thredds_creator = "DOD/USAF/SMC > Space and Missile Systems Center (SMC), U.S. Air Force, U.S. Department of Defense";
 :thredds_contributor = "DOC/NOAA/NESDIS/NGDC > National Geophysical Data Center, NESDIS, NOAA, U.S. Department of Commerce";
 :thredds_contributor_role = "archive";
 :thredds_publisher = "DOC/NOAA/NESDIS/NGDC > National Geophysical Data Center, NESDIS, NOAA, U.S. Department of Commerce";
 :thredds_publisher_url = "http://dmsp.ngdc.noaa.gov/";
 :thredds_publisher_email = "ngdc.dmsp@noaa.gov";
 :thredds_summary = "This dataset contains data from the DMSP F14 satellite OLS instrument and includes both visible smooth and thermal smooth imagery with 2.7km resolution. The start time for this data is 2003-07-19T22:30:31.371GMT and the northerly equatorial crossing longitude is 320.54.  The DMSP satellite is a polar-orbiting satellite crossing the equator, depending on the satellite, at either dawn/dusk or noon/midnight. This data is in the NOAA/NGDC DMSP archive format.";
 :thredds_history = "";
 :thredds_timeCoverage_start = "2003-07-19T22:30:31.371GMT";
 :thredds_timeCoverage_end = "2003-07-19T22:35:21.836GMT";
 :thredds_geospatialCoverage = "Polar orbit with northerly equatorial crossing at longitude 320.55.";
}