netcdf dods://localhost:8082/dts/test.02 {
  variables:
    ubyte b(25);

    int i32(25);

    uint ui32(25);

    short i16(25);

    ushort ui16(25);

    float f32(25);

    double f64(25);

    String s(25);

    String u(25);

}
