netcdf dods://iridl.ldeo.columbia.edu/SOURCES/.NOAA/.NCEP/.CPC/.GLOBAL/.daily/dods {
 dimensions:
   nmiss = 7;
   time = 13791;
   lon = 144;
   lat = 73;
 variables:
   float nmiss(nmiss=7);
     :pointwidth = 1.0f; // float
     :gridtype = 0; // int
     :units = "unitless";
   float time(time=13791);
     :calendar = "standard";
     :pointwidth = 1.0f; // float
     :gridtype = 0; // int
     :units = "days since 1974-01-01";
   float lon(lon=144);
     :long_name = "Longitude";
     :actual_range = 0.0f, 360.0f; // float
     :pointwidth = 2.5f; // float
     :modulus = 360.0f; // float
     :standard_name = "longitude";
     :axis = "X";
     :gridtype = 1; // int
     :units = "degree_east";
   float lat(lat=73);
     :axis = "Y";
     :long_name = "Latitude";
     :standard_name = "latitude";
     :pointwidth = 2.5f; // float
     :actual_range = 90.0f, -90.0f; // float
     :gridtype = 0; // int
     :units = "degree_north";
   short info(time=13791, nmiss=7);
     :_CoordinateAxes = "time nmiss ";
     :valid_range = 0, 10512; // int
     :units = "unitless";
     :missing_value = 32766S; // short
     :long_name = "Missing";
   short olr(time=13791, lat=73, lon=144);
     :_CoordinateAxes = "time lat lon ";
     :var_desc = "Outgoing Longwave Radiation";
     :scale_factor = 0.01f; // float
     :actual_range = 98.5f, 315.0f; // float
     :dataset = "NOAA Interpolated OLR";
     :units = "W/m2";
     :unpacked_valid_range = 0.0f, 500.0f; // float
     :valid_range = -32765, 17235; // int
     :level_desc = "Other";
     :statistic = "Mean";
     :precision = 2; // int
     :add_offset = 327.65f; // float
     :missing_value = 32766S; // short
     :long_name = "Daily OLR";
     :parent_stat = "Individual Obs";

 :Conventions = "COARDS";
 :NCO = "4.0.0";
 :history = "Tue May 10 11:37:33 2005: ncatted -a missing_value,info,o,s,32766 /Datasets/interp_OLR/olr.day.mean.nc", "/home/hoop/crdc/oldCRDC2COARDSv3/oldCRDC2COARDS Sat Dec  9 01:36:34 1995 from olr.7494.nc", "created 08/24/94 by C. Smith (netCDF2.3)";
 :description = "Data is interpolated in time and space from NOAA twice-daily OLR values and averaged to once daily";
 :platform = "Observation";
 :title = "Daily Mean Interpolated OLR";
 :reference = "Liebmann and Smith (Bulletin of the American Meteorological Society 1996)";
 :references = "Liebmann_Smith1996";
 :dataset_documentation.html = "http://iridl.ldeo.columbia.edu/SOURCES/.NOAA/.NCEP/.CPC/.GLOBAL/.daily/.dataset_documentation.html";
}
