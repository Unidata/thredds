netcdf test_misc1 {
dimensions:
	lat = 6 ;
	lon = 4 ;
	time = UNLIMITED ; // (0 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
	double time(time) ;
		time:units = "seconds since 2009-01-01" ;
	float pr(time, lat, lon) ;
		pr:standard_name = "air_pressure_at_sea_level" ;
		pr:units = "hPa" ;

// global attributes:
		:title = "example for workshop" ;
}
