netcdf dods://iridl.ldeo.columbia.edu/SOURCES/.NOAA/.NCEP/.CPC/.GLOBAL/.daily/dods {
 dimensions:
   nmiss = 7;
   time = 14063;
   lon = 144;
   lat = 73;
 variables:
   float nmiss(nmiss=7);
     :pointwidth = 1.0f; // float
     :gridtype = 0; // int
     :units = "unitless";
   float time(time=14063);
     :calendar = "standard";
     :pointwidth = 1.0f; // float
     :gridtype = 0; // int
     :units = "days since 1974-01-01";
   float lon(lon=144);
     :standard_name = "longitude";
     :modulus = 360.0f; // float
     :pointwidth = 2.5f; // float
     :axis = "X";
     :actual_range = 0.0f, 360.0f; // float
     :long_name = "Longitude";
     :gridtype = 1; // int
     :units = "degree_east";
   float lat(lat=73);
     :standard_name = "latitude";
     :actual_range = 90.0f, -90.0f; // float
     :long_name = "Latitude";
     :axis = "Y";
     :pointwidth = 2.5f; // float
     :gridtype = 0; // int
     :units = "degree_north";
   short info(time=14063, nmiss=7);
     :_CoordinateAxes = "time nmiss ";
     :units = "unitless";
     :missing_value = 32766S; // short
     :long_name = "Missing";
     :valid_range = 0, 10512; // int
   short olr(time=14063, lat=73, lon=144);
     :_CoordinateAxes = "time lat lon ";
     :valid_range = -32765, 17235; // int
     :long_name = "Daily OLR";
     :level_desc = "Other";
     :dataset = "NOAA Interpolated OLR";
     :units = "W/m2";
     :scale_factor = 0.01f; // float
     :statistic = "Mean";
     :precision = 2; // int
     :var_desc = "Outgoing Longwave Radiation";
     :parent_stat = "Individual Obs";
     :actual_range = 94.625f, 316.5f; // float
     :add_offset = 327.65f; // float
     :missing_value = 32766S; // short
     :unpacked_valid_range = 0.0f, 500.0f; // float
 // global attributes:
 :reference = "Liebmann and Smith (Bulletin of the American Meteorological Society 1996)";
 :references = "Liebmann_Smith1996";
 :dataset_documentation.html = "http://iridl.ldeo.columbia.edu/SOURCES/.NOAA/.NCEP/.CPC/.GLOBAL/.daily/.dataset_documentation.html";
 :NCO = "4.0.0";
 :history = "Tue May 10 11:37:33 2005: ncatted -a missing_value,info,o,s,32766 /Datasets/interp_OLR/olr.day.mean.nc", "/home/hoop/crdc/oldCRDC2COARDSv3/oldCRDC2COARDS Sat Dec  9 01:36:34 1995 from olr.7494.nc", "created 08/24/94 by C. Smith (netCDF2.3)";
 :platform = "Observation";
 :title = "Daily Mean Interpolated OLR";
 :description = "Data is interpolated in time and space from NOAA twice-daily OLR values and averaged to once daily";
 :Conventions = "COARDS";
}
