netcdf dods://remotetest.unidata.ucar.edu/dts/test.22?exp.ThreeD[5:1:7][5:8][1:3] {
  dimensions:
    x = 3;
    y = 4;
    z = 3;
  variables:

    Structure {
      double x(x=3);
      double y(y=4);
      double z(z=3);
      double ThreeD(x=3, y=4, z=3);
        :_CoordinateAxes = "x y z ";
    } exp;


}
