netcdf test_vlen4 {
types:
  int(*) v_t ;
  compound c_t {
    v_t f1(2) ;
  }; // c_t
variables:
	c_t v1 ;
data:

 v1 = {{{1, 3, 5, 7}, {100, 200}}} ;
}
