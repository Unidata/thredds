netcdf dods://remotetest.unidata.ucar.edu/thredds/dodsC/testdods/K1VHR.nc {
 dimensions:
   GeoX = 4;
   time = 1;
   GeoY = 4;
 variables:
   int GeoX(GeoX=4);
     :long_name = "x-coordinate in Cartesian system";
     :axis = "X";

   float time(time=1);
     :units = "hours since 2000-01-01 00:00:00";

   int GeoY(GeoY=4);
     :long_name = "y-coordinate in Cartesian system";
     :axis = "Y";


 group: Science_Data {

   group: Geolocation_Information {
     variables:
       short Latitude(GeoY=4, GeoX=4);
         :_CoordinateAxes = "GeoY GeoX ";
         :scale_factor = 0.01f; // float
         :units = "degrees_north";
         :_FillValue = 32767S; // short
         :standard_name = "latitude";
         :add_offset = 0.0f; // float
         :_ChunkSize = 1400, 1400; // int
       short Longitude(GeoY=4, GeoX=4);
         :_CoordinateAxes = "GeoY GeoX ";
         :_FillValue = 32767S; // short
         :scale_factor = 0.01f; // float
         :units = "degrees_east";
         :add_offset = 0.0f; // float
         :standard_name = "longitude";
         :_ChunkSize = 1400, 1400; // int
   }

   group: Geophysical_Parameter {
     variables:
       float OLR(time=1, GeoY=4, GeoX=4);
         :_CoordinateAxes = "time GeoY GeoX ";
         :coordinates = "time Latitude Longitude";
         :long_name = "Outgoing Longwave Radiation";
         :standard_name = "Outgoing Longwave Radiation";
         :_FillValue = -999.0f; // float
         :units = "W.m-2";
         :_ChunkSize = 1, 936, 1400; // int
   }
 }
 // global attributes:
 :institute = "Space Applications Center, ISRO";
 :source = "Very High Resolution Radiometer (VHRR)";
 :conventions = "CF-1.6";
 :title = "K1VHR_05JUL2012_0700_L2B";
 :Product_Metadata47Unique_Id = "K1VHR_05JUL2012_0700";
 :Product_Metadata47Product_Creation_Time = "2012-07-08T13:05:32";
 :Product_Metadata47Output_Format = "hdf5-1.8.8";
 :Product_Metadata47HDF_Product_File_Name = "K1VHR_05JUL2012_0700_L2B_OLR.h5";
 :Product_Metadata47Station_Id = "BES";
 :Product_Metadata47Ground_Station = "BES,SAC/ISRO,Ahmedabad,INDIA.";
 :Product_Metadata47Servo_Correction = "X";
 :Product_Metadata47Detector_Normalization = "Y";
 :Product_Metadata47Shear_Correction = "X";
 :Product_Metadata47Inoperable_Detectors = "Y";
 :Product_Metadata47Dropped_Lines = "Y";
 :Product_Metadata47EW_Count_Variation = "X";
 :Product_Metadata47Product_Type = "GEOPHY";
 :Product_Metadata47Sensor_Id = "VHR";
 :Product_Metadata47Sensor_Name = "VHRR";
 :Product_Metadata47Acquisition_Date = "05JUL2012";
 :Product_Metadata47Acquisition_Time_in_GMT = "0700";
 :Product_Metadata47Processing_Level = "L2B";
 :Product_Metadata47Satellite_Name = "KALPANA-1";
 :Product_Metadata47Location_of_Satellite(degrees) = 74.0f; // float
 :Product_Metadata47Imaging_Mode = "NORMAL FRAME";
 :Product_Metadata47Nominal_Altitude(km) = 36000.0f; // float
 :Product_Metadata47Predicted_Altitude(km) = 35793.98f; // float
 :Product_Metadata47Black_Body_Strategy_Used_for_Thermal_IR_Band = "Current Black Body Line";
 :Product_Metadata47Nominal_Pixel_Stepping_Angle(degrees) = 0.012707; // double
 :Product_Metadata47Pixel_Stepping_Angle(degrees) = 0.012707; // double
 :Product_Metadata47Nominal_Line_Stepping_Angle(degrees) = 0.012784; // double
 :Product_Metadata47Line_Stepping_Angle(degrees) = 0.012784; // double
 :Product_Metadata47Field_of_View(degrees) = 19.82292; // double
 :Product_Metadata47Nominal_Central_Point_Coordinates(degrees)_Latitude_Longitude = 0.0, 74.0; // double
 :Product_Metadata47Predicted_Central_Point_Coordinates(degrees)_Latitude_Longitude = 1.726647, 73.899302; // double
}
