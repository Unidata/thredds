netcdf group.test2 {
 group: g1 {
   variables:
     int i32;
 }
 group: g2 {
   variables:
     int i32;
 }
}
