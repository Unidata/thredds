netcdf testgrid2 {
dimensions:
  time = 2;
variables:
  double var(time,time) ;
  float time(time);
data:
  var = 0.0, 1.0, 2.0, 3.0, 4.0;
  time = 17.0, 23.0;
}
